localparam IDLE = 2'b00;
localparam HAZARD = 2'b01;
localparam TURN = 2'b10;

localparam LEFT = 0;
localparam RIGHT = 1;
