localparam IDLE = 2'b00;
localparam HAZARD = 2'b01;
localparam LTURN = 2'b10;
localparam RTURN = 2'b11;

localparam LEFT = 0;
localparam RIGHT = 1;
