localparam IDLE = 2'b00;
localparam HAZARD = 2'b01;
localparam TURN = 2'b10;
