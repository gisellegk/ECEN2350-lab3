module blinker(input clock, input state, output [2:0]LEDs);

endmodule